module sprite(
	input clk,
	input reset,

	input red_in,
	input green_in,
	input blue_in,

	output red_out,
	output green_out,
	output blue_out
);

endmodule
